`timescale 1 ns/1 ns
module Sdcontroller_tb;

reg clk, reset;

// Instantiate UUT
SDcontroller UUT(


endmodule;